//--------------------------------------------------------------------------------------------------------
// Module  : command_processor
// Function: receive 8 bytes from AXI-stream slave, then take various actions
//--------------------------------------------------------------------------------------------------------

module command_processor (
	input  wire        rstn,
	input  wire        clk,
	// AXI-stream slave
	output wire        i_tready,
	input  wire        i_tvalid,
	input  wire [ 7:0] i_tdata,
	// AXI-stream master
	input  wire        o_tready,
	output wire        o_tvalid,
	output wire [31:0] o_tdata,
	output wire [ 3:0] o_tkeep,
	output wire        o_tlast,
	 
	output reg pllreset,
	 
	output reg [7:0]	spitx,
	input  reg [7:0]	spirx,
	input  reg 			spitxready,
	output reg			spitxdv,
	input  reg			spirxdv,
	output reg [7:0]	spics, // which chip to talk to
	
	input wire			locked, // clock is locked
	
	input wire [139:0] lvds1bits, lvds2bits, lvds3bits, lvds4bits,// rx_in[0] drives data to rx_out[(J-1)..0], rx_in[1] drives data to the next J number of bits on rx_out
	input wire			clklvds, // clk1, runs at LVDS bit rate (ADC clk input rate) / 2
	output reg			lvds1wr,
	output reg			lvds1rd,
	input wire			lvds1wrfull,
	input wire			lvds1wrempty,
	input wire			lvds1rdfull,
	input wire			lvds1rdempty,
	output reg [559:0] lvds1bitsfifoout, //output bits to fifo
	input wire [559:0] lvds1bitsfifoin, // input bits from fifo
	input wire [19:0] lvdsbits_o2, lvdsbits_other,
	
	output reg[2:0] phasecounterselect, // Dynamic phase shift counter Select. 000:all 001:M 010:C0 011:C1 100:C2 101:C3 110:C4. Registered in the rising edge of scanclk.
	output reg phaseupdown=1, // Dynamic phase shift direction; 1:UP, 0:DOWN. Registered in the PLL on the rising edge of scanclk.
	output reg [3:0] phasestep,
	output reg scanclk=0,

	output reg [2:0] spimisossel=0, //which spimiso to listen to
	output reg [11:0]	debugout,  // for debugging
	input wire [3:0]	overrange,  //ORA0,A1,B0,B1
	
	output reg [1:0] spi_mode=0,
	
	input wire [7:0] boardin,
	output wire [7:0] boardout,
	output reg spireset_L,
	input wire clk50, // needed while doing pllreset,
	input wire lvdsin_trig,
	output reg lvdsout_trig=0,
	output reg clkswitch=0,
	input wire lvdsin_spare[2],
	output reg lvdsout_spare[2]
);

integer version = 14; // firmware version

assign debugout[0] = locked;
assign debugout[1] = spics[4];
assign debugout[2] = spics[5];
assign debugout[3] = phaseupdown;
assign debugout[4] = overrange[0];
assign debugout[5] = overrange[1];
assign debugout[6] = overrange[2];
assign debugout[7] = overrange[3];
assign debugout[11:8] = state;

assign lvdsout_trig = lvdsin_trig;

//for clock phase
reg[7:0] pllclock_counter=0;
reg[7:0] scanclk_cycles=0;
  

//variables in clk domain
localparam [3:0] INIT=4'd0, RX=4'd1, PROCESS=4'd2, TX_DATA_CONST=4'd3, TX_DATA1=4'd4, TX_DATA2=4'd5, TX_DATA3=4'd6, TX_DATA4=4'd7, PLLCLOCK=4'd8;
reg [ 3:0]	state = INIT;
reg [ 3:0]	rx_counter = 0;
reg [ 7:0]	rx_data[7:0];
integer		length = 0;
reg [ 3:0]	spistate = 0;
reg [5:0]	channel = 0;
reg [3:0]	spicscounter = 0;

//variables in clklvds domain
reg [ 2:0]  acqstate=0;
reg [15:0]	triggercounter=0, triggercounter_sync=0;
reg [15:0]	eventcounter=0, eventcounter_sync=0;
reg [15:0]	lengthtotake=0, lengthtotake_sync=0;
reg 			triggerlive=0, triggerlive_sync=0;
reg			didreadout=0, didreadout_sync=0;
reg [ 7:0]	triggertype=0, triggertype_sync=0;
reg signed [11:0]  lowerthresh=-12'd10, upperthresh=12'd10;

reg signed [11:0]  samplevalue[40];
reg [1:0] sampleclkstr[40];

integer i;
always @ (posedge clklvds) begin
	
	triggerlive_sync <= triggerlive;
	lengthtotake_sync <= lengthtotake;
	triggertype_sync <= triggertype;
	didreadout_sync <= didreadout;

	for (i=0;i<10;i=i+1) begin
		samplevalue[i]  <= {lvds1bits[110+i],lvds1bits[100+i],lvds1bits[90+i],lvds1bits[80+i],lvds1bits[70+i],lvds1bits[60+i],lvds1bits[50+i],lvds1bits[40+i],lvds1bits[30+i],lvds1bits[20+i],lvds1bits[10+i],lvds1bits[0+i]};
		sampleclkstr[i] <= {lvds1bits[130+i],lvds1bits[120+i]};
		samplevalue[10+i]  <= {lvds2bits[110+i],lvds2bits[100+i],lvds2bits[90+i],lvds2bits[80+i],lvdsbits_other[0+i],lvdsbits_other[10+i],lvds2bits[50+i],lvds2bits[40+i],lvds2bits[30+i],lvds2bits[20+i],lvds2bits[10+i],lvds2bits[0+i]};
		sampleclkstr[10+i] <= {lvds2bits[130+i],lvds2bits[120+i]};
		samplevalue[20+i]  <= {lvds3bits[110+i],lvds3bits[100+i],lvds3bits[90+i],lvds3bits[80+i],lvds3bits[70+i],lvds3bits[60+i],lvds3bits[50+i],lvds3bits[40+i],lvds3bits[30+i],lvds3bits[20+i],lvds3bits[10+i],lvds3bits[0+i]};
		sampleclkstr[20+i] <= {lvds3bits[130+i],lvds3bits[120+i]};
		samplevalue[30+i]  <= {lvdsbits_o2[0+i],lvds4bits[100+i],lvds4bits[90+i],lvds4bits[80+i],lvds4bits[70+i],lvds4bits[60+i],lvds4bits[50+i],lvds4bits[40+i],lvds4bits[30+i],lvds4bits[20+i],lvds4bits[10+i],lvds4bits[0+i]};
		sampleclkstr[30+i] <= {lvds4bits[130+i],lvds4bits[120+i]};
	end
end

always @ (posedge clklvds or negedge rstn)
 if (~rstn) begin
	lvds1wr <= 1'b0;
	acqstate <= 3'd0;
 end else begin
	case (acqstate)
	0 : begin // ready
		lvds1wr <= 1'b0;
		triggercounter<=0;
		if (triggerlive_sync) begin
			if (triggertype_sync==8'd1) acqstate <= 3'd1; // threshold trigger
			else acqstate <= 3'd3; // go straight to taking data, no trigger, triggertype==0
		end
	end
	1 : begin // ready for first part of trigger condition to be met
		if (samplevalue[0]<lowerthresh) acqstate <= 3'd2;
	end
	2 : begin // ready for second part of trigger condition to be met
		if (samplevalue[0]>upperthresh) acqstate <= 3'd3;
	end
	3 : begin // taking data
		lvds1bitsfifoout <= {
		sampleclkstr[39],samplevalue[39],sampleclkstr[38],samplevalue[38],sampleclkstr[37],samplevalue[37],sampleclkstr[36],samplevalue[36],sampleclkstr[35],samplevalue[35],sampleclkstr[34],samplevalue[34],sampleclkstr[33],samplevalue[33],sampleclkstr[32],samplevalue[32],sampleclkstr[31],samplevalue[31],sampleclkstr[30],samplevalue[30],
		sampleclkstr[29],samplevalue[29],sampleclkstr[28],samplevalue[28],sampleclkstr[27],samplevalue[27],sampleclkstr[26],samplevalue[26],sampleclkstr[25],samplevalue[25],sampleclkstr[24],samplevalue[24],sampleclkstr[23],samplevalue[23],sampleclkstr[22],samplevalue[22],sampleclkstr[21],samplevalue[21],sampleclkstr[20],samplevalue[20],
		sampleclkstr[19],samplevalue[19],sampleclkstr[18],samplevalue[18],sampleclkstr[17],samplevalue[17],sampleclkstr[16],samplevalue[16],sampleclkstr[15],samplevalue[15],sampleclkstr[14],samplevalue[14],sampleclkstr[13],samplevalue[13],sampleclkstr[12],samplevalue[12],sampleclkstr[11],samplevalue[11],sampleclkstr[10],samplevalue[10],	
		sampleclkstr[9],samplevalue[9],sampleclkstr[8],samplevalue[8],sampleclkstr[7],samplevalue[7],sampleclkstr[6],samplevalue[6],sampleclkstr[5],samplevalue[5],sampleclkstr[4],samplevalue[4],sampleclkstr[3],samplevalue[3],sampleclkstr[2],samplevalue[2],sampleclkstr[1],samplevalue[1],sampleclkstr[0],samplevalue[0]
		};
		//lvds1bitsfifoout <= {56{triggercounter[9:0]}}; // for testing the queue
		if ((!lvds1wrfull) && triggercounter<lengthtotake_sync) begin
			lvds1wr <= 1'b1;
			triggercounter<=triggercounter+16'd1;
		end
		else begin
			lvds1wr <= 1'b0;
			eventcounter <= eventcounter+16'd1;
			acqstate <= 3'd4;
		end
	end
	4 : begin // ready to be read out
		triggercounter<= -16'd1;
		if (didreadout_sync) acqstate <= 3'd0;
	end
	default : begin
		acqstate <= 3'd0;
	end
	endcase
 end
 
integer overrange_counter[4];
always @ (posedge clk) begin
	
	triggercounter_sync <= triggercounter;
	eventcounter_sync <= eventcounter;
	
	if (overrange[0]) overrange_counter[0]<=overrange_counter[0]+1;
	if (overrange[1]) overrange_counter[1]<=overrange_counter[1]+1;
	if (overrange[2]) overrange_counter[2]<=overrange_counter[2]+1;
	if (overrange[3]) overrange_counter[3]<=overrange_counter[3]+1;
end

reg [1:0] pllresetstate=0;
reg pllreset2=0;
always @ (posedge clk50) begin
	case (pllresetstate)
   0 : begin
		if (pllreset2) begin
			pllreset<=1'b1;
			pllresetstate<=2'd1;
		end
	end
	1 : begin
		pllreset<=1'b0;
		if (!pllreset2) pllresetstate<=2'd0;
	end
	endcase
end

always @ (posedge clk or negedge rstn)
 if (~rstn) begin
	state  <= INIT;
 end else begin
 
  case (state)
   INIT : begin
		spireset_L <= 1'b1;
		pllreset2 <= 1'b0;
		lvds1rd <= 1'b0;
   	rx_counter <= 0;
		length <= 0;
		spistate <= 0;
		spitxdv <= 1'b0;
		spics <= 8'hff;
		channel <= 6'd0;
		triggerlive <= 1'b0;
		didreadout <= 1'b0;
		state <= RX;
	end
  
	RX : if (i_tvalid) begin // get 8 bytes
		rx_data[rx_counter] <= i_tdata;
		if (rx_counter==7) begin
			 state <= PROCESS;
			 rx_counter <= 0;
		end
		else rx_counter <= rx_counter+4'd1;
	end
	
	PROCESS : begin // do something, based on the command in the first byte
		case (rx_data[0])
			
		0 : begin // send a length of bytes
			didreadout <= 1'b1; // tell it we have read out this event
			length <= {rx_data[7],rx_data[6],rx_data[5],rx_data[4]};
			state <= TX_DATA1;
		end
		
		1 : begin // sets length of data to take, activates trigger for new event if we don't alrady have one
			triggertype <= rx_data[1]; // while we're at it, set the trigger type
			lengthtotake <= {rx_data[5],rx_data[4]};
			if (triggercounter_sync == 0) triggerlive <= 1'b1; // gets reset in INIT state
			//else triggerlive <= 1'b0;
			o_tdata <= {eventcounter_sync,triggercounter_sync}; // return triggercounter, so we can see if we have an event ready to be read out
			length <= 4;
			o_tvalid <= 1'b1;
			state <= TX_DATA_CONST;
		end
		
		2 : begin // reads version or other info
			if (rx_data[1]==0) o_tdata <= version;
			if (rx_data[1]==1) o_tdata <= {boardin,boardin,boardin,boardin};
			if (rx_data[1]==2) o_tdata <= overrange_counter[rx_data[2][1:0]];
			length <= 4;
			o_tvalid <= 1'b1;
			state <= TX_DATA_CONST;
		end
		
		3 : begin // SPI command
			case (spistate)			
			0 : begin
				spimisossel <= rx_data[1][2:0]; // select requested data from chip
				spics[rx_data[1][2:0]]<=1'b0; //select requested chip
				spitx <= rx_data[2];//first byte to send
				
				if (spicscounter==4'd5) begin // wait a bit for cs to go low
					spicscounter<=4'd0;
					spistate <= 4'd1;
				end
				else spicscounter<=spicscounter+4'd1;
			end
			1 : begin
				if (spitxready) begin
					spitxdv <= 1'b1;
					if (rx_data[7]==2) spistate <= 4'd4; //sending 2 bytes
					else spistate <= 4'd2; // sending more than 2 bytes
				end
			end
			2 : begin
				spitxdv <= 1'b0;
				spitx <= rx_data[3];//second byte to send
				spistate <= 4'd3;
			end
			3 : begin
				if (spitxready) begin
					spitxdv <= 1'b1;
					spistate <= 4'd4;
				end
			end
			4 : begin
				spitxdv <= 1'b0;
				spitx <= rx_data[4];//third byte to send (ignored during read)
				spistate <= 4'd5;
			end
			5 : begin
				if (spitxready) begin
					spitxdv <= 1'b1;
					if (rx_data[7]==4) spistate <= 4'd6; // send the 4th byte
					else spistate <= 4'd8; // skip the 4th byte
				end
			end
			6 : begin
				spitxdv <= 1'b0;
				spitx <= rx_data[5];//fourth byte to send
				spistate <= 4'd7;
			end
			7 : begin
				if (spitxready) begin
					spitxdv <= 1'b1;
					spistate <= 4'd8;
				end
			end
			8 : begin
				spitxdv <= 1'b0;
				if (spirxdv) begin
					spistate <= 4'd9;
					o_tdata <= spirx; // send back the SPI data read
				end
			end
			9 : begin
				if (spicscounter==4'd15) begin // wait a bit before setting cs high
					spicscounter<=4'd0;
					spistate <= 4'd0;
					length <= 4;
					o_tvalid <= 1'b1;
					state <= TX_DATA_CONST;		
				end
				else spicscounter<=spicscounter+4'd1;
			end
			default : spistate <= 4'd0;
			endcase
		end
		
		4 : begin // set SPI_MODE (see SPI_Master.v)
			spireset_L <= 1'b0;
			spi_mode <= rx_data[1][1:0];
			o_tdata <= rx_data[1];
			length <= 4;
			o_tvalid <= 1'b1;
			state <= TX_DATA_CONST;
		end
		
		5 : begin // reset plls
			pllreset2 <= 1'b1;
			o_tdata <= 33;
			length <= 4;
			o_tvalid <= 1'b1;
			state <= TX_DATA_CONST;
		end
		
		6 : begin
			phasecounterselect<=rx_data[2][2:0];// 000:all 001:M 010:C0 011:C1 100:C2 101:C3 110:C4. 
			phaseupdown<=rx_data[3][0]; // up or down
			scanclk<=1'b0; // start low
			phasestep[rx_data[1]]<=1'b1; // assert!
			pllclock_counter<=0;
			scanclk_cycles<=0;
			state<=PLLCLOCK;
		end
		
		7 : begin // try to switch clocks
			clkswitch <= ~clkswitch;
			o_tdata <= {8'd0,8'd0,8'd0,7'd0,~clkswitch};
			length <= 4;
			o_tvalid <= 1'b1;
			state <= TX_DATA_CONST;
		end
		
		default: // some command we didn't know
			state <= RX;
			
		endcase
	end
	
	TX_DATA_CONST : if (o_tready) begin
		if (length >= 4) begin
			length <= length - 16'd4;
		end else begin
			length <= 0;
			o_tvalid <= 1'b0;
			state <= INIT;
		end
	end
	
	TX_DATA1 : begin //channel==0
		o_tvalid <= 1'b0;
		if (o_tready) begin
			if (lvds1rdempty) begin // wait for data
				lvds1rd <= 1'b0;
			end
			else begin
				lvds1rd <= 1'b1;
				state <= TX_DATA2;
			end
		end
	end
	
	TX_DATA2 : begin // wait for read
		lvds1rd <= 1'b0;
		o_tvalid <= 1'b0;
		if (o_tready) begin
			state <= TX_DATA3;
		end
	end
	
	TX_DATA3 : begin
		lvds1rd <= 1'b0;
		if (o_tready) begin
			o_tvalid <= 1'b1;
			if (channel==48) o_tdata <= {16'hbeef,16'hdead};//marker
			else if (channel==46) o_tdata  <= {
				12'd0,
				lvds1bitsfifoin[14*39+12 +: 2], //sampleclkstr39
				lvds1bitsfifoin[14*38+12 +: 2],lvds1bitsfifoin[14*37+12 +: 2],lvds1bitsfifoin[14*36+12 +: 2],lvds1bitsfifoin[14*35+12 +: 2],lvds1bitsfifoin[14*34+12 +: 2],lvds1bitsfifoin[14*33+12 +: 2],lvds1bitsfifoin[14*32+12 +: 2],lvds1bitsfifoin[14*31+12 +: 2],
				lvds1bitsfifoin[14*30+12 +: 2], //sampleclkstr30
				};
			else if (channel==44) o_tdata  <= {
				12'd0,
				lvds1bitsfifoin[14*29+12 +: 2], //sampleclkstr29
				lvds1bitsfifoin[14*28+12 +: 2],lvds1bitsfifoin[14*27+12 +: 2],lvds1bitsfifoin[14*26+12 +: 2],lvds1bitsfifoin[14*25+12 +: 2],lvds1bitsfifoin[14*24+12 +: 2],lvds1bitsfifoin[14*23+12 +: 2],lvds1bitsfifoin[14*22+12 +: 2],lvds1bitsfifoin[14*21+12 +: 2],
				lvds1bitsfifoin[14*20+12 +: 2], //sampleclkstr20
				};
			else if (channel==42) o_tdata  <= {
				12'd0,
				lvds1bitsfifoin[14*19+12 +: 2], //sampleclkstr19
				lvds1bitsfifoin[14*18+12 +: 2],lvds1bitsfifoin[14*17+12 +: 2],lvds1bitsfifoin[14*16+12 +: 2],lvds1bitsfifoin[14*15+12 +: 2],lvds1bitsfifoin[14*14+12 +: 2],lvds1bitsfifoin[14*13+12 +: 2],lvds1bitsfifoin[14*12+12 +: 2],lvds1bitsfifoin[14*11+12 +: 2],
				lvds1bitsfifoin[14*10+12 +: 2], //sampleclkstr10
				};
			else if (channel==40) o_tdata  <= {
				12'd0,
				lvds1bitsfifoin[14*9+12 +: 2], //sampleclkstr9
				lvds1bitsfifoin[14*8+12 +: 2],lvds1bitsfifoin[14*7+12 +: 2],lvds1bitsfifoin[14*6+12 +: 2],lvds1bitsfifoin[14*5+12 +: 2],lvds1bitsfifoin[14*4+12 +: 2],lvds1bitsfifoin[14*3+12 +: 2],lvds1bitsfifoin[14*2+12 +: 2],lvds1bitsfifoin[14*1+12 +: 2],
				lvds1bitsfifoin[14*0+12 +: 2], //sampleclkstr0
				};
			else o_tdata  <= {4'd0, lvds1bitsfifoin[14*(channel+1) +: 12], 4'd0, lvds1bitsfifoin[14*channel +: 12]};
			channel<=channel+6'd2;
			state <= TX_DATA4;
		end
	end
	
	TX_DATA4 : begin
		lvds1rd <= 1'b0;
		if (o_tready) begin
			o_tvalid <= 1'b0;
			if (length >= 4) begin
				length <= length - 16'd4;
				if (channel==50) begin
					channel <= 0;
					state <= TX_DATA1;
				end
				else state <= TX_DATA3;
			end 
			else begin
				length <= 0;
				channel<=0;
				state <= RX;
			end
		end
	end
	
	PLLCLOCK : begin // to step the clock phase, you have to toggle scanclk a few times
		pllclock_counter <= pllclock_counter+8'd1;
		if (pllclock_counter[4]) begin
			scanclk <= ~scanclk;
			pllclock_counter <= 0;
			scanclk_cycles <= scanclk_cycles+8'd1;
			if (scanclk_cycles>5) phasestep[rx_data[1]] <= 1'b0; // deassert!
			if (scanclk_cycles>7) state <= INIT;
		end
	end
	
	default :
		state <= RX;
	
  endcase
 end

assign i_tready = (state == RX);
assign o_tkeep  = (length>=4) ? 4'b1111 :
                  (length==3) ? 4'b0111 :
                  (length==2) ? 4'b0011 :
                  (length==1) ? 4'b0001 :
                 /*length==0*/  4'b0000;
assign o_tlast  = (length>=4) ? 1'b0 : 1'b1;
endmodule
